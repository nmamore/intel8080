/*
* @file intel8080_top.sv
* @brief top-level file for the Intel 8080
* @author Nicholas Amore namore7@gmail.com
* @date Created 1/2/2023
*/

`timescale 1ns / 100ps

module intel8080_top
(
    input logic clk50M_i,
    input logic rst_ni
    
);

endmodule